//============================================================================
//
//  AUTHOR      : YoungBeom Kim
//  SPEC        :
//  HISTORY     : 2023-11-08 오전 12:13:28
//
//      Copyright (c) 2023 Crypto Optimization & Application LAb. MIT license
//
//============================================================================


//Problem : Implement the wire following circuit:

module top_module
(
	input	in	,
		
	output	out
);

assign	out = in;

endmodule