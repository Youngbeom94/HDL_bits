//============================================================================
//
//  AUTHOR      : YoungBeom Kim
//  SPEC        :
//  HISTORY     : 2024-10-01 오후 7:16:06
//
//      Copyright (c) 2024 Crypto & Security Engineering Laboratory. MIT license
//
//============================================================================

// synthesis verilog_input_version verilog_2001
module top_module 
( 
    input		[2:0] sel	, 
    input		[3:0] data0	,
    input		[3:0] data1	,
    input		[3:0] data2	,
    input		[3:0] data3	,
    input		[3:0] data4	,
    input		[3:0] data5	,
    output	reg [3:0] out   
);//

wire [3:0] imm;

assign	imm =	sel == 3'b000 ? data0 : 
				sel == 3'b001 ? data1 : 
				sel == 3'b010 ? data2 : 
				sel == 3'b011 ? data3 : 
				sel == 3'b100 ? data4 : 
				sel == 3'b101 ? data5 : 0;				

	// Another Solution
    always@(*) begin  
        out <= imm;
    end
    
//    basic solution => This is a combinational circuit
//    always@(*) begin  
//        case(sel)
//        	3'b000:	out <= data0;
//        	3'b001:	out <= data1;
//        	3'b010:	out <= data2;
//        	3'b011:	out <= data3;
//        	3'b100:	out <= data4;
//        	3'b101:	out <= data5;
//        	default:out <= 0;        	
//    	endcase
//    end

endmodule