//============================================================================
//
//  AUTHOR      : YoungBeom Kim
//  SPEC        :
//  HISTORY     : 2024-06-12 오후 5:52:00
//
//      Copyright (c) 2024 Crypto & Security Engineering Laboratory. MIT license
//
//============================================================================


// Problem
// Solution
module top_module
(
	input		a	,
	input		b	,
	input		c	,
	output		w	,
	output		x	,
	output		y	,
	output		z	
);                                                                                                      

	assign w = a;
	assign x = b;
	assign y = b;	
	assign z = c;	
       
endmodule

// Anothor solution provied by HDL_bits.