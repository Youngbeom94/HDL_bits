//============================================================================
//
//  AUTHOR      : YoungBeom Kim
//  SPEC        :
//  HISTORY     : 2023-11-08 오전 12:55:50
//
//      Copyright (c) 2023 Crypto Optimization & Application LAb. MIT license
//
//============================================================================


//Problem : Create a 4-bit wide, 256-to-1 multiplexer. The 256 4-bit inputs are all packed into a single 1024-bit input vector. sel=0 should select bits in[3:0], sel=1 selects bits in[7:4], sel=2 selects bits in[11:8], etc.
// My solution
module top_module
(
	input	[1023:0]	in	,
	input	[7:0]		sel	,
		
	output	[3:0]		out	
);                                                                                                      

assign	out = (sel == 0  ) ? in[4*(0  +1)-1:4*0  ] : (sel == 1  ) ? in[4*(1  +1)-1:4*1  ] : (sel == 2  ) ? in[4*(2  +1)-1:4*2  ] : (sel == 3  ) ? in[4*(3  +1)-1:4*3  ] : 
              (sel == 4  ) ? in[4*(4  +1)-1:4*4  ] : (sel == 5  ) ? in[4*(5  +1)-1:4*5  ] : (sel == 6  ) ? in[4*(6  +1)-1:4*6  ] : (sel == 7  ) ? in[4*(7  +1)-1:4*7  ] : 
              (sel == 8  ) ? in[4*(8  +1)-1:4*8  ] : (sel == 9  ) ? in[4*(9  +1)-1:4*9  ] : (sel == 10 ) ? in[4*(10 +1)-1:4*10 ] : (sel == 11 ) ? in[4*(11 +1)-1:4*11 ] : 
              (sel == 12 ) ? in[4*(12 +1)-1:4*12 ] : (sel == 13 ) ? in[4*(13 +1)-1:4*13 ] : (sel == 14 ) ? in[4*(14 +1)-1:4*14 ] : (sel == 15 ) ? in[4*(15 +1)-1:4*15 ] : 
              (sel == 16 ) ? in[4*(16 +1)-1:4*16 ] : (sel == 17 ) ? in[4*(17 +1)-1:4*17 ] : (sel == 18 ) ? in[4*(18 +1)-1:4*18 ] : (sel == 19 ) ? in[4*(19 +1)-1:4*19 ] : 
              (sel == 20 ) ? in[4*(20 +1)-1:4*20 ] : (sel == 21 ) ? in[4*(21 +1)-1:4*21 ] : (sel == 22 ) ? in[4*(22 +1)-1:4*22 ] : (sel == 23 ) ? in[4*(23 +1)-1:4*23 ] : 
              (sel == 24 ) ? in[4*(24 +1)-1:4*24 ] : (sel == 25 ) ? in[4*(25 +1)-1:4*25 ] : (sel == 26 ) ? in[4*(26 +1)-1:4*26 ] : (sel == 27 ) ? in[4*(27 +1)-1:4*27 ] : 
              (sel == 28 ) ? in[4*(28 +1)-1:4*28 ] : (sel == 29 ) ? in[4*(29 +1)-1:4*29 ] : (sel == 30 ) ? in[4*(30 +1)-1:4*30 ] : (sel == 31 ) ? in[4*(31 +1)-1:4*31 ] : 
              (sel == 32 ) ? in[4*(32 +1)-1:4*32 ] : (sel == 33 ) ? in[4*(33 +1)-1:4*33 ] : (sel == 34 ) ? in[4*(34 +1)-1:4*34 ] : (sel == 35 ) ? in[4*(35 +1)-1:4*35 ] : 
              (sel == 36 ) ? in[4*(36 +1)-1:4*36 ] : (sel == 37 ) ? in[4*(37 +1)-1:4*37 ] : (sel == 38 ) ? in[4*(38 +1)-1:4*38 ] : (sel == 39 ) ? in[4*(39 +1)-1:4*39 ] : 
              (sel == 40 ) ? in[4*(40 +1)-1:4*40 ] : (sel == 41 ) ? in[4*(41 +1)-1:4*41 ] : (sel == 42 ) ? in[4*(42 +1)-1:4*42 ] : (sel == 43 ) ? in[4*(43 +1)-1:4*43 ] : 
              (sel == 44 ) ? in[4*(44 +1)-1:4*44 ] : (sel == 45 ) ? in[4*(45 +1)-1:4*45 ] : (sel == 46 ) ? in[4*(46 +1)-1:4*46 ] : (sel == 47 ) ? in[4*(47 +1)-1:4*47 ] : 
              (sel == 48 ) ? in[4*(48 +1)-1:4*48 ] : (sel == 49 ) ? in[4*(49 +1)-1:4*49 ] : (sel == 50 ) ? in[4*(50 +1)-1:4*50 ] : (sel == 51 ) ? in[4*(51 +1)-1:4*51 ] : 
              (sel == 52 ) ? in[4*(52 +1)-1:4*52 ] : (sel == 53 ) ? in[4*(53 +1)-1:4*53 ] : (sel == 54 ) ? in[4*(54 +1)-1:4*54 ] : (sel == 55 ) ? in[4*(55 +1)-1:4*55 ] : 
              (sel == 56 ) ? in[4*(56 +1)-1:4*56 ] : (sel == 57 ) ? in[4*(57 +1)-1:4*57 ] : (sel == 58 ) ? in[4*(58 +1)-1:4*58 ] : (sel == 59 ) ? in[4*(59 +1)-1:4*59 ] : 
              (sel == 60 ) ? in[4*(60 +1)-1:4*60 ] : (sel == 61 ) ? in[4*(61 +1)-1:4*61 ] : (sel == 62 ) ? in[4*(62 +1)-1:4*62 ] : (sel == 63 ) ? in[4*(63 +1)-1:4*63 ] : 
              (sel == 64 ) ? in[4*(64 +1)-1:4*64 ] : (sel == 65 ) ? in[4*(65 +1)-1:4*65 ] : (sel == 66 ) ? in[4*(66 +1)-1:4*66 ] : (sel == 67 ) ? in[4*(67 +1)-1:4*67 ] : 
              (sel == 68 ) ? in[4*(68 +1)-1:4*68 ] : (sel == 69 ) ? in[4*(69 +1)-1:4*69 ] : (sel == 70 ) ? in[4*(70 +1)-1:4*70 ] : (sel == 71 ) ? in[4*(71 +1)-1:4*71 ] : 
              (sel == 72 ) ? in[4*(72 +1)-1:4*72 ] : (sel == 73 ) ? in[4*(73 +1)-1:4*73 ] : (sel == 74 ) ? in[4*(74 +1)-1:4*74 ] : (sel == 75 ) ? in[4*(75 +1)-1:4*75 ] : 
              (sel == 76 ) ? in[4*(76 +1)-1:4*76 ] : (sel == 77 ) ? in[4*(77 +1)-1:4*77 ] : (sel == 78 ) ? in[4*(78 +1)-1:4*78 ] : (sel == 79 ) ? in[4*(79 +1)-1:4*79 ] : 
              (sel == 80 ) ? in[4*(80 +1)-1:4*80 ] : (sel == 81 ) ? in[4*(81 +1)-1:4*81 ] : (sel == 82 ) ? in[4*(82 +1)-1:4*82 ] : (sel == 83 ) ? in[4*(83 +1)-1:4*83 ] : 
              (sel == 84 ) ? in[4*(84 +1)-1:4*84 ] : (sel == 85 ) ? in[4*(85 +1)-1:4*85 ] : (sel == 86 ) ? in[4*(86 +1)-1:4*86 ] : (sel == 87 ) ? in[4*(87 +1)-1:4*87 ] : 
              (sel == 88 ) ? in[4*(88 +1)-1:4*88 ] : (sel == 89 ) ? in[4*(89 +1)-1:4*89 ] : (sel == 90 ) ? in[4*(90 +1)-1:4*90 ] : (sel == 91 ) ? in[4*(91 +1)-1:4*91 ] : 
              (sel == 92 ) ? in[4*(92 +1)-1:4*92 ] : (sel == 93 ) ? in[4*(93 +1)-1:4*93 ] : (sel == 94 ) ? in[4*(94 +1)-1:4*94 ] : (sel == 95 ) ? in[4*(95 +1)-1:4*95 ] : 
              (sel == 96 ) ? in[4*(96 +1)-1:4*96 ] : (sel == 97 ) ? in[4*(97 +1)-1:4*97 ] : (sel == 98 ) ? in[4*(98 +1)-1:4*98 ] : (sel == 99 ) ? in[4*(99 +1)-1:4*99 ] : 
              (sel == 100) ? in[4*(100+1)-1:4*100] : (sel == 101) ? in[4*(101+1)-1:4*101] : (sel == 102) ? in[4*(102+1)-1:4*102] : (sel == 103) ? in[4*(103+1)-1:4*103] : 
              (sel == 104) ? in[4*(104+1)-1:4*104] : (sel == 105) ? in[4*(105+1)-1:4*105] : (sel == 106) ? in[4*(106+1)-1:4*106] : (sel == 107) ? in[4*(107+1)-1:4*107] : 
              (sel == 108) ? in[4*(108+1)-1:4*108] : (sel == 109) ? in[4*(109+1)-1:4*109] : (sel == 110) ? in[4*(110+1)-1:4*110] : (sel == 111) ? in[4*(111+1)-1:4*111] : 
              (sel == 112) ? in[4*(112+1)-1:4*112] : (sel == 113) ? in[4*(113+1)-1:4*113] : (sel == 114) ? in[4*(114+1)-1:4*114] : (sel == 115) ? in[4*(115+1)-1:4*115] : 
              (sel == 116) ? in[4*(116+1)-1:4*116] : (sel == 117) ? in[4*(117+1)-1:4*117] : (sel == 118) ? in[4*(118+1)-1:4*118] : (sel == 119) ? in[4*(119+1)-1:4*119] : 
              (sel == 120) ? in[4*(120+1)-1:4*120] : (sel == 121) ? in[4*(121+1)-1:4*121] : (sel == 122) ? in[4*(122+1)-1:4*122] : (sel == 123) ? in[4*(123+1)-1:4*123] : 
              (sel == 124) ? in[4*(124+1)-1:4*124] : (sel == 125) ? in[4*(125+1)-1:4*125] : (sel == 126) ? in[4*(126+1)-1:4*126] : (sel == 127) ? in[4*(127+1)-1:4*127] : 
              (sel == 128) ? in[4*(128+1)-1:4*128] : (sel == 129) ? in[4*(129+1)-1:4*129] : (sel == 130) ? in[4*(130+1)-1:4*130] : (sel == 131) ? in[4*(131+1)-1:4*131] : 
              (sel == 132) ? in[4*(132+1)-1:4*132] : (sel == 133) ? in[4*(133+1)-1:4*133] : (sel == 134) ? in[4*(134+1)-1:4*134] : (sel == 135) ? in[4*(135+1)-1:4*135] : 
              (sel == 136) ? in[4*(136+1)-1:4*136] : (sel == 137) ? in[4*(137+1)-1:4*137] : (sel == 138) ? in[4*(138+1)-1:4*138] : (sel == 139) ? in[4*(139+1)-1:4*139] : 
              (sel == 140) ? in[4*(140+1)-1:4*140] : (sel == 141) ? in[4*(141+1)-1:4*141] : (sel == 142) ? in[4*(142+1)-1:4*142] : (sel == 143) ? in[4*(143+1)-1:4*143] : 
              (sel == 144) ? in[4*(144+1)-1:4*144] : (sel == 145) ? in[4*(145+1)-1:4*145] : (sel == 146) ? in[4*(146+1)-1:4*146] : (sel == 147) ? in[4*(147+1)-1:4*147] : 
              (sel == 148) ? in[4*(148+1)-1:4*148] : (sel == 149) ? in[4*(149+1)-1:4*149] : (sel == 150) ? in[4*(150+1)-1:4*150] : (sel == 151) ? in[4*(151+1)-1:4*151] : 
              (sel == 152) ? in[4*(152+1)-1:4*152] : (sel == 153) ? in[4*(153+1)-1:4*153] : (sel == 154) ? in[4*(154+1)-1:4*154] : (sel == 155) ? in[4*(155+1)-1:4*155] : 
              (sel == 156) ? in[4*(156+1)-1:4*156] : (sel == 157) ? in[4*(157+1)-1:4*157] : (sel == 158) ? in[4*(158+1)-1:4*158] : (sel == 159) ? in[4*(159+1)-1:4*159] : 
              (sel == 160) ? in[4*(160+1)-1:4*160] : (sel == 161) ? in[4*(161+1)-1:4*161] : (sel == 162) ? in[4*(162+1)-1:4*162] : (sel == 163) ? in[4*(163+1)-1:4*163] : 
              (sel == 164) ? in[4*(164+1)-1:4*164] : (sel == 165) ? in[4*(165+1)-1:4*165] : (sel == 166) ? in[4*(166+1)-1:4*166] : (sel == 167) ? in[4*(167+1)-1:4*167] : 
              (sel == 168) ? in[4*(168+1)-1:4*168] : (sel == 169) ? in[4*(169+1)-1:4*169] : (sel == 170) ? in[4*(170+1)-1:4*170] : (sel == 171) ? in[4*(171+1)-1:4*171] : 
              (sel == 172) ? in[4*(172+1)-1:4*172] : (sel == 173) ? in[4*(173+1)-1:4*173] : (sel == 174) ? in[4*(174+1)-1:4*174] : (sel == 175) ? in[4*(175+1)-1:4*175] : 
              (sel == 176) ? in[4*(176+1)-1:4*176] : (sel == 177) ? in[4*(177+1)-1:4*177] : (sel == 178) ? in[4*(178+1)-1:4*178] : (sel == 179) ? in[4*(179+1)-1:4*179] : 
              (sel == 180) ? in[4*(180+1)-1:4*180] : (sel == 181) ? in[4*(181+1)-1:4*181] : (sel == 182) ? in[4*(182+1)-1:4*182] : (sel == 183) ? in[4*(183+1)-1:4*183] : 
              (sel == 184) ? in[4*(184+1)-1:4*184] : (sel == 185) ? in[4*(185+1)-1:4*185] : (sel == 186) ? in[4*(186+1)-1:4*186] : (sel == 187) ? in[4*(187+1)-1:4*187] : 
              (sel == 188) ? in[4*(188+1)-1:4*188] : (sel == 189) ? in[4*(189+1)-1:4*189] : (sel == 190) ? in[4*(190+1)-1:4*190] : (sel == 191) ? in[4*(191+1)-1:4*191] : 
              (sel == 192) ? in[4*(192+1)-1:4*192] : (sel == 193) ? in[4*(193+1)-1:4*193] : (sel == 194) ? in[4*(194+1)-1:4*194] : (sel == 195) ? in[4*(195+1)-1:4*195] : 
              (sel == 196) ? in[4*(196+1)-1:4*196] : (sel == 197) ? in[4*(197+1)-1:4*197] : (sel == 198) ? in[4*(198+1)-1:4*198] : (sel == 199) ? in[4*(199+1)-1:4*199] : 
              (sel == 200) ? in[4*(200+1)-1:4*200] : (sel == 201) ? in[4*(201+1)-1:4*201] : (sel == 202) ? in[4*(202+1)-1:4*202] : (sel == 203) ? in[4*(203+1)-1:4*203] : 
              (sel == 204) ? in[4*(204+1)-1:4*204] : (sel == 205) ? in[4*(205+1)-1:4*205] : (sel == 206) ? in[4*(206+1)-1:4*206] : (sel == 207) ? in[4*(207+1)-1:4*207] : 
              (sel == 208) ? in[4*(208+1)-1:4*208] : (sel == 209) ? in[4*(209+1)-1:4*209] : (sel == 210) ? in[4*(210+1)-1:4*210] : (sel == 211) ? in[4*(211+1)-1:4*211] : 
              (sel == 212) ? in[4*(212+1)-1:4*212] : (sel == 213) ? in[4*(213+1)-1:4*213] : (sel == 214) ? in[4*(214+1)-1:4*214] : (sel == 215) ? in[4*(215+1)-1:4*215] : 
              (sel == 216) ? in[4*(216+1)-1:4*216] : (sel == 217) ? in[4*(217+1)-1:4*217] : (sel == 218) ? in[4*(218+1)-1:4*218] : (sel == 219) ? in[4*(219+1)-1:4*219] : 
              (sel == 220) ? in[4*(220+1)-1:4*220] : (sel == 221) ? in[4*(221+1)-1:4*221] : (sel == 222) ? in[4*(222+1)-1:4*222] : (sel == 223) ? in[4*(223+1)-1:4*223] : 
              (sel == 224) ? in[4*(224+1)-1:4*224] : (sel == 225) ? in[4*(225+1)-1:4*225] : (sel == 226) ? in[4*(226+1)-1:4*226] : (sel == 227) ? in[4*(227+1)-1:4*227] : 
              (sel == 228) ? in[4*(228+1)-1:4*228] : (sel == 229) ? in[4*(229+1)-1:4*229] : (sel == 230) ? in[4*(230+1)-1:4*230] : (sel == 231) ? in[4*(231+1)-1:4*231] : 
              (sel == 232) ? in[4*(232+1)-1:4*232] : (sel == 233) ? in[4*(233+1)-1:4*233] : (sel == 234) ? in[4*(234+1)-1:4*234] : (sel == 235) ? in[4*(235+1)-1:4*235] : 
              (sel == 236) ? in[4*(236+1)-1:4*236] : (sel == 237) ? in[4*(237+1)-1:4*237] : (sel == 238) ? in[4*(238+1)-1:4*238] : (sel == 239) ? in[4*(239+1)-1:4*239] : 
              (sel == 240) ? in[4*(240+1)-1:4*240] : (sel == 241) ? in[4*(241+1)-1:4*241] : (sel == 242) ? in[4*(242+1)-1:4*242] : (sel == 243) ? in[4*(243+1)-1:4*243] : 
              (sel == 244) ? in[4*(244+1)-1:4*244] : (sel == 245) ? in[4*(245+1)-1:4*245] : (sel == 246) ? in[4*(246+1)-1:4*246] : (sel == 247) ? in[4*(247+1)-1:4*247] : 
              (sel == 248) ? in[4*(248+1)-1:4*248] : (sel == 249) ? in[4*(249+1)-1:4*249] : (sel == 250) ? in[4*(250+1)-1:4*250] : (sel == 251) ? in[4*(251+1)-1:4*251] : 
              (sel == 252) ? in[4*(252+1)-1:4*252] : (sel == 253) ? in[4*(253+1)-1:4*253] : (sel == 254) ? in[4*(254+1)-1:4*254] : (sel == 255) ? in[4*(255+1)-1:4*255] : 'b0;
       
endmodule

// Anothor solution provied by HDL_bits.
module top_module
(
	input	[1023:0]	in	,
	input	[7:0]		sel	,
		
	output	[3:0]		out	
);   

	// We can't part-select multiple bits without an error, but we can select one bit at a time,
	// four times, then concatenate them together.
	assign out = {in[sel*4+3], in[sel*4+2], in[sel*4+1], in[sel*4+0]};

	// Alternatively, "indexed vector part select" works better, but has an unfamiliar syntax:
	// assign out = in[sel*4 +: 4];		// Select starting at index "sel*4", then select a total width of 4 bits with increasing (+:) index number.
	// assign out = in[sel*4+3 -: 4];	// Select starting at index "sel*4+3", then select a total width of 4 bits with decreasing (-:) index number.
	// Note: The width (4 in this case) must be constant.

endmodule