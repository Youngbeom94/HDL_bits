//============================================================================
//
//  AUTHOR      : YoungBeom Kim
//  SPEC        :
//  HISTORY     : 2024-10-01 오후 7:02:57
//
//      Copyright (c) 2024 Crypto & Security Engineering Laboratory. MIT license
//
//============================================================================

// synthesis verilog_input_version verilog_2001
module top_module 
(
    input      cpu_overheated,
    output reg shut_off_computer,
    
    input      arrived,
    input      gas_tank_empty,
    output reg keep_driving 
);

    always @(*) begin
        if (cpu_overheated) begin
           shut_off_computer <= 1;
        end
        else begin
        	shut_off_computer <= 0;
    	end
    end

    always @(*) begin
        if (~arrived) begin
           keep_driving = ~gas_tank_empty;
        end
        else begin
        	keep_driving = 0;
    	end
    end

endmodule