//============================================================================
//
//  AUTHOR      : YoungBeom Kim
//  SPEC        :
//  HISTORY     : 2024-06-12 오후 5:44:28
//
//      Copyright (c) 2024 Crypto & Security Engineering Laboratory. MIT license
//
//============================================================================


// Problem
// Solution
module top_module
(
	input		in	,			
	output		out	
);                                                                                                      

	assign out = in;
       
endmodule

// Anothor solution provied by HDL_bits.